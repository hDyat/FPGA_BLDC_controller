module rpm_lut (
	datain,
	dataout
);
	
	input [7:0] datain;
	output reg [9:0] dataout;

	always @ (datain)
		case(datain)
			8'd0:	dataout = 10'd0;
			8'd1: dataout = 10'd4;
			8'd2: dataout = 10'd8;
			8'd3: dataout = 10'd12;
			8'd4: dataout = 10'd16;
			8'd5: dataout = 10'd20;
			8'd6: dataout = 10'd24;
			8'd7: dataout = 10'd28;
			8'd8: dataout = 10'd32;
			8'd9: dataout = 10'd36;
			8'd10: dataout = 10'd40;
			8'd11: dataout = 10'd44;
			8'd12: dataout = 10'd48;
			8'd13: dataout = 10'd52;
			8'd14: dataout = 10'd56;
			8'd15: dataout = 10'd60;
			8'd16: dataout = 10'd64;
			8'd17: dataout = 10'd68;
			8'd18: dataout = 10'd72;
			8'd19: dataout = 10'd76;
			8'd20: dataout = 10'd80;
			8'd21: dataout = 10'd84;
			8'd22: dataout = 10'd88;
			8'd23: dataout = 10'd92;
			8'd24: dataout = 10'd96;
			8'd25: dataout = 10'd100;
			8'd26: dataout = 10'd104;
			8'd27: dataout = 10'd108;
			8'd28: dataout = 10'd112;
			8'd29: dataout = 10'd116;
			8'd30: dataout = 10'd120;
			8'd31: dataout = 10'd124;
			8'd32: dataout = 10'd128;
			8'd33: dataout = 10'd132;
			8'd34: dataout = 10'd136;
			8'd35: dataout = 10'd140;
			8'd36: dataout = 10'd144;
			8'd37: dataout = 10'd148;
			8'd38: dataout = 10'd152;
			8'd39: dataout = 10'd156;
			8'd40: dataout = 10'd160;
			8'd41: dataout = 10'd164;
			8'd42: dataout = 10'd168;
			8'd43: dataout = 10'd172;
			8'd44: dataout = 10'd176;
			8'd45: dataout = 10'd180;
			8'd46: dataout = 10'd184;
			8'd47: dataout = 10'd188;
			8'd48: dataout = 10'd192;
			8'd49: dataout = 10'd196;
			8'd50: dataout = 10'd200;
			8'd51: dataout = 10'd204;
			8'd52: dataout = 10'd208;
			8'd53: dataout = 10'd212;
			8'd54: dataout = 10'd216;
			8'd55: dataout = 10'd220;
			8'd56: dataout = 10'd224;
			8'd57: dataout = 10'd228;
			8'd58: dataout = 10'd232;
			8'd59: dataout = 10'd236;
			8'd60: dataout = 10'd240;
			8'd61: dataout = 10'd244;
			8'd62: dataout = 10'd248;
			8'd63: dataout = 10'd252;
			8'd64: dataout = 10'd256;
			8'd65: dataout = 10'd260;
			8'd66: dataout = 10'd264;
			8'd67: dataout = 10'd268;
			8'd68: dataout = 10'd272;
			8'd69: dataout = 10'd276;
			8'd70: dataout = 10'd280;
			8'd71: dataout = 10'd284;
			8'd72: dataout = 10'd288;
			8'd73: dataout = 10'd292;
			8'd74: dataout = 10'd296;
			8'd75: dataout = 10'd300;
			8'd76: dataout = 10'd304;
			8'd77: dataout = 10'd308;
			8'd78: dataout = 10'd312;
			8'd79: dataout = 10'd316;
			8'd80: dataout = 10'd320;
			8'd81: dataout = 10'd324;
			8'd82: dataout = 10'd328;
			8'd83: dataout = 10'd332;
			8'd84: dataout = 10'd336;
			8'd85: dataout = 10'd340;
			8'd86: dataout = 10'd344;
			8'd87: dataout = 10'd348;
			8'd88: dataout = 10'd352;
			8'd89: dataout = 10'd356;
			8'd90: dataout = 10'd360;
			8'd91: dataout = 10'd364;
			8'd92: dataout = 10'd368;
			8'd93: dataout = 10'd372;
			8'd94: dataout = 10'd376;
			8'd95: dataout = 10'd380;
			8'd96: dataout = 10'd384;
			8'd97: dataout = 10'd388;
			8'd98: dataout = 10'd392;
			8'd99: dataout = 10'd396;
			8'd100: dataout = 10'd400;
			8'd101: dataout = 10'd404;
			8'd102: dataout = 10'd408;
			8'd103: dataout = 10'd412;
			8'd104: dataout = 10'd416;
			8'd105: dataout = 10'd420;
			8'd106: dataout = 10'd424;
			8'd107: dataout = 10'd428;
			8'd108: dataout = 10'd432;
			8'd109: dataout = 10'd436;
			8'd110: dataout = 10'd440;
			8'd111: dataout = 10'd444;
			8'd112: dataout = 10'd448;
			8'd113: dataout = 10'd452;
			8'd114: dataout = 10'd456;
			8'd115: dataout = 10'd460;
			8'd116: dataout = 10'd464;
			8'd117: dataout = 10'd468;
			8'd118: dataout = 10'd472;
			8'd119: dataout = 10'd476;
			8'd120: dataout = 10'd480;
			8'd121: dataout = 10'd484;
			8'd122: dataout = 10'd488;
			8'd123: dataout = 10'd491;
			8'd124: dataout = 10'd496;
			8'd125: dataout = 10'd500;
			8'd126: dataout = 10'd504;
			8'd127: dataout = 10'd508;
			8'd128: dataout = 10'd512;
			8'd129: dataout = 10'd516;
			8'd130: dataout = 10'd520;
			8'd131: dataout = 10'd524;
			8'd132: dataout = 10'd528;
			8'd133: dataout = 10'd532;
			8'd134: dataout = 10'd536;
			8'd135: dataout = 10'd540;
			8'd136: dataout = 10'd544;
			8'd137: dataout = 10'd548;
			8'd138: dataout = 10'd552;
			8'd139: dataout = 10'd556;
			8'd140: dataout = 10'd560;
			8'd141: dataout = 10'd564;
			8'd142: dataout = 10'd568;
			8'd143: dataout = 10'd572;
			8'd144: dataout = 10'd576;
			8'd145: dataout = 10'd580;
			8'd146: dataout = 10'd584;
			8'd147: dataout = 10'd588;
			8'd148: dataout = 10'd592;
			8'd149: dataout = 10'd596;
			8'd150: dataout = 10'd600;
			8'd151: dataout = 10'd604;
			8'd152: dataout = 10'd608;
			8'd153: dataout = 10'd612;
			8'd154: dataout = 10'd616;
			8'd155: dataout = 10'd620;
			8'd156: dataout = 10'd624;
			8'd157: dataout = 10'd628;
			8'd158: dataout = 10'd632;
			8'd159: dataout = 10'd636;
			8'd160: dataout = 10'd640;
			8'd161: dataout = 10'd644;
			8'd162: dataout = 10'd648;
			8'd163: dataout = 10'd652;
			8'd164: dataout = 10'd656;
			8'd165: dataout = 10'd660;
			8'd166: dataout = 10'd664;
			8'd167: dataout = 10'd668;
			8'd168: dataout = 10'd672;
			8'd169: dataout = 10'd676;
			8'd170: dataout = 10'd680;
			8'd171: dataout = 10'd684;
			8'd172: dataout = 10'd688;
			8'd173: dataout = 10'd692;
			8'd174: dataout = 10'd696;
			8'd175: dataout = 10'd700;
			8'd176: dataout = 10'd704;
			8'd177: dataout = 10'd708;
			8'd178: dataout = 10'd712;
			8'd179: dataout = 10'd716;
			8'd180: dataout = 10'd720;
			8'd181: dataout = 10'd724;
			8'd182: dataout = 10'd728;
			8'd183: dataout = 10'd732;
			8'd184: dataout = 10'd736;
			8'd185: dataout = 10'd740;
			8'd186: dataout = 10'd744;
			8'd187: dataout = 10'd748;
			8'd188: dataout = 10'd752;
			8'd189: dataout = 10'd756;
			8'd190: dataout = 10'd760;
			8'd191: dataout = 10'd764;
			8'd192: dataout = 10'd768;
			8'd193: dataout = 10'd772;
			8'd194: dataout = 10'd776;
			8'd195: dataout = 10'd780;
			8'd196: dataout = 10'd784;
			8'd197: dataout = 10'd788;
			8'd198: dataout = 10'd792;
			8'd199: dataout = 10'd796;
			8'd200: dataout = 10'd800;
			default: ;
		endcase
endmodule
