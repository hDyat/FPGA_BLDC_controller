module rpm_lut (D, Q);
    input      [10:0] D;
    output reg [10:0] Q;

    always @ (D)
        case(D)
            11'h0:	Q = 11'h0;
            11'h1:	Q = 11'ha;
            11'h2:	Q = 11'h14;
            11'h3:	Q = 11'h1e;
            11'h4:	Q = 11'h28;
            11'h5:	Q = 11'h32;
            11'h6:	Q = 11'h3c;
            11'h7:	Q = 11'h46;
            11'h8:	Q = 11'h50;
            11'h9:	Q = 11'h5a;
            11'ha:	Q = 11'h64;
            11'hb:	Q = 11'h6e;
            11'hc:	Q = 11'h78;
            11'hd:	Q = 11'h82;
            11'he:	Q = 11'h8c;
            11'hf:	Q = 11'h96;
            11'h10:	Q = 11'ha0;
            11'h11:	Q = 11'haa;
            11'h12:	Q = 11'hb4;
            11'h13:	Q = 11'hbe;
            11'h14:	Q = 11'hc8;
            11'h15:	Q = 11'hd2;
            11'h16:	Q = 11'hdc;
            11'h17:	Q = 11'he6;
            11'h18:	Q = 11'hf0;
            11'h19:	Q = 11'hfa;
            11'h1a:	Q = 11'h104;
            11'h1b:	Q = 11'h10e;
            11'h1c:	Q = 11'h118;
            11'h1d:	Q = 11'h122;
            11'h1e:	Q = 11'h12c;
            11'h1f:	Q = 11'h136;
            11'h20:	Q = 11'h140;
            11'h21:	Q = 11'h14a;
            11'h22:	Q = 11'h154;
            11'h23:	Q = 11'h15e;
            11'h24:	Q = 11'h168;
            11'h25:	Q = 11'h172;
            11'h26:	Q = 11'h17c;
            11'h27:	Q = 11'h186;
            11'h28:	Q = 11'h190;
            11'h29:	Q = 11'h19a;
            11'h2a:	Q = 11'h1a4;
            11'h2b:	Q = 11'h1ae;
            11'h2c:	Q = 11'h1b8;
            11'h2d:	Q = 11'h1c2;
            11'h2e:	Q = 11'h1cc;
            11'h2f:	Q = 11'h1d6;
            11'h30:	Q = 11'h1e0;
            11'h31:	Q = 11'h1ea;
            11'h32:	Q = 11'h1f4;
            11'h33:	Q = 11'h1fe;
            11'h34:	Q = 11'h208;
            11'h35:	Q = 11'h212;
            11'h36:	Q = 11'h21c;
            11'h37:	Q = 11'h226;
            11'h38:	Q = 11'h230;
            11'h39:	Q = 11'h23a;
            11'h3a:	Q = 11'h244;
            11'h3b:	Q = 11'h24e;
            11'h3c:	Q = 11'h258;
            11'h3d:	Q = 11'h262;
            11'h3e:	Q = 11'h26c;
            11'h3f:	Q = 11'h276;
            11'h40:	Q = 11'h280;
            11'h41:	Q = 11'h28a;
            11'h42:	Q = 11'h294;
            11'h43:	Q = 11'h29e;
            11'h44:	Q = 11'h2a8;
            11'h45:	Q = 11'h2b2;
            11'h46:	Q = 11'h2bc;
            11'h47:	Q = 11'h2c6;
            11'h48:	Q = 11'h2d0;
            11'h49:	Q = 11'h2da;
            11'h4a:	Q = 11'h2e4;
            11'h4b:	Q = 11'h2ee;
            11'h4c:	Q = 11'h2f8;
            11'h4d:	Q = 11'h302;
            11'h4e:	Q = 11'h30c;
            11'h4f:	Q = 11'h316;
            11'h50:	Q = 11'h320;
            11'h51:	Q = 11'h32a;
            11'h52:	Q = 11'h334;
            11'h53:	Q = 11'h33e;
            11'h54:	Q = 11'h348;
            11'h55:	Q = 11'h352;
            11'h56:	Q = 11'h35c;
            11'h57:	Q = 11'h366;
            11'h58:	Q = 11'h370;
            11'h59:	Q = 11'h37a;
            11'h5a:	Q = 11'h384;
            11'h5b:	Q = 11'h38e;
            11'h5c:	Q = 11'h398;
            11'h5d:	Q = 11'h3a2;
            11'h5e:	Q = 11'h3ac;
            11'h5f:	Q = 11'h3b6;
            11'h60:	Q = 11'h3c0;
            11'h61:	Q = 11'h3ca;
            11'h62:	Q = 11'h3d4;
            11'h63:	Q = 11'h3de;
            11'h64:	Q = 11'h3e8;
            11'h65:	Q = 11'h3f2;
            11'h66:	Q = 11'h3fc;
            11'h67:	Q = 11'h406;
            11'h68:	Q = 11'h410;
            11'h69:	Q = 11'h41a;
            11'h6a:	Q = 11'h424;
            11'h6b:	Q = 11'h42e;
            11'h6c:	Q = 11'h438;
            11'h6d:	Q = 11'h442;
            11'h6e:	Q = 11'h44c;
            11'h6f:	Q = 11'h456;
            11'h70:	Q = 11'h460;
            11'h71:	Q = 11'h46a;
            11'h72:	Q = 11'h474;
            11'h73:	Q = 11'h47e;
            11'h74:	Q = 11'h488;
            11'h75:	Q = 11'h492;
            11'h76:	Q = 11'h49c;
            11'h77:	Q = 11'h4a6;
            11'h78:	Q = 11'h4b0;
            11'h79:	Q = 11'h4ba;
            11'h7a:	Q = 11'h4c4;
            11'h7b:	Q = 11'h4ce;
            11'h7c:	Q = 11'h4d8;
            11'h7d:	Q = 11'h4e2;
            11'h7e:	Q = 11'h4ec;
            11'h7f:	Q = 11'h4f6;
            11'h80:	Q = 11'h500;
            11'h81:	Q = 11'h50a;
            11'h82:	Q = 11'h514;
            11'h83:	Q = 11'h51e;
            11'h84:	Q = 11'h528;
            11'h85:	Q = 11'h532;
            11'h86:	Q = 11'h53c;
            11'h87:	Q = 11'h546;
            11'h88:	Q = 11'h550;
            11'h89:	Q = 11'h55a;
            11'h8a:	Q = 11'h564;
            11'h8b:	Q = 11'h56e;
            11'h8c:	Q = 11'h578;
            11'h8d:	Q = 11'h582;
            11'h8e:	Q = 11'h58c;
            11'h8f:	Q = 11'h596;
            11'h90:	Q = 11'h5a0;
            11'h91:	Q = 11'h5aa;
            11'h92:	Q = 11'h5b4;
            11'h93:	Q = 11'h5be;
            11'h94:	Q = 11'h5c8;
            11'h95:	Q = 11'h5d2;
            11'h96:	Q = 11'h5dc;
            11'h97:	Q = 11'h5e6;
            11'h98:	Q = 11'h5f0;
            11'h99:	Q = 11'h5fa;
            11'h9a:	Q = 11'h604;
            11'h9b:	Q = 11'h60e;
            11'h9c:	Q = 11'h618;
            11'h9d:	Q = 11'h622;
            11'h9e:	Q = 11'h62c;
            11'h9f:	Q = 11'h636;
            11'ha0:	Q = 11'h640;
            11'ha1:	Q = 11'h64a;
            11'ha2:	Q = 11'h654;
            11'ha3:	Q = 11'h65e;
            11'ha4:	Q = 11'h668;
            11'ha5:	Q = 11'h672;
            11'ha6:	Q = 11'h67c;
            11'ha7:	Q = 11'h686;
            11'ha8:	Q = 11'h690;
            11'ha9:	Q = 11'h69a;
            11'haa:	Q = 11'h6a4;
            11'hab:	Q = 11'h6ae;
            11'hac:	Q = 11'h6b8;
            11'had:	Q = 11'h6c2;
            11'hae:	Q = 11'h6cc;
            11'haf:	Q = 11'h6d6;
            11'hb0:	Q = 11'h6e0;
            11'hb1:	Q = 11'h6ea;
            11'hb2:	Q = 11'h6f4;
            11'hb3:	Q = 11'h6fe;
            11'hb4:	Q = 11'h708;
            11'hb5:	Q = 11'h712;
            11'hb6:	Q = 11'h71c;
            11'hb7:	Q = 11'h726;
            11'hb8:	Q = 11'h730;
            11'hb9:	Q = 11'h73a;
            11'hba:	Q = 11'h744;
            11'hbb:	Q = 11'h74e;
            11'hbc:	Q = 11'h758;
            11'hbd:	Q = 11'h762;
            11'hbe:	Q = 11'h76c;
            11'hbf:	Q = 11'h776;
            11'hc0:	Q = 11'h780;
            11'hc1:	Q = 11'h78a;
            11'hc2:	Q = 11'h794;
            11'hc3:	Q = 11'h79e;
            11'hc4:	Q = 11'h7a8;
            11'hc5:	Q = 11'h7b2;
            11'hc6:	Q = 11'h7bc;
            11'hc7:	Q = 11'h7c6;
            11'hc8:	Q = 11'h7d0;
            default:	Q = 11'hxxx;
        endcase
endmodule
