module unipolar_pwm (
	
);

endmodule